-------------------------------------------------------------------------------
--
-- Title       : ALU
-- Design      : ALU
-- Author      : C3C John Paul Terragnoli 
-- Company     : usafa
--
-------------------------------------------------------------------------------
--
-- File        : ALU.vhd
-- Generated   : Apr 7 11:16:54 2041
-- From        : interface description file
--
-------------------------------------------------------------------------------
--
-- Description : Holds the logic for the ALU. 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {ALU} architecture {ALU}}

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ALU is
	 port(
		 OpSel : in STD_LOGIC_VECTOR(2 downto 0);
		 Data : in STD_LOGIC_VECTOR(3 downto 0);
		 Accumulator : in STD_LOGIC_VECTOR(3 downto 0);
		 Result : out STD_LOGIC_VECTOR(3 downto 0)
	     );
end ALU;

--}} End of automatically maintained section

architecture ALU of ALU is	   


begin
	
-- fill in details to create result as a function of Data and Accumulator, based on OpSel.
 -- e.g : Build a multiplexer choosing between the eight ALU operations.  Either use a case statement (and thus a process)
 --       or a conditional signal assignment statement ( x <= Y when <condition> else . . .)
 -- ALU Operations are defined as:
 -- OpSel : Function
--  0     : AND
--  1     : NEG (2s complement)
--  2     : NOT (invert)
--  3     : ROR
--  4     : OR
--  5     : IN
--  6     : ADD
--  7     : LD
--aluswitch: process (Accumulator, Data, OpSel)
--        begin
--		  -- enter your if/then/else or case statements here
--		end process;

-- OR, enter your conditional signal statement here
Result <= (Data and Accumulator) when (Opsel = "000") else
			((not Accumulator)+ "001") when (Opsel =  "001") else
			(not Accumulator) when (Opsel = "010") else
			--this one will be awesome if it works.  
			(accumulator(0)&accumulator(3) &accumulator(2)&accumulator(1)) when (Opsel = "011") else
			(Data or Accumulator) when (Opsel  = "100") else
			(Data) when (Opsel = "101") else
			(Data + Accumulator) when (Opsel = "110") else
			(Data) when (Opsel = "111") else
			--nothing specified, put what is in the accumulator in the result.  
			Accumulator; 	
end ALU;

